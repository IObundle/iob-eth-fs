// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UUT_DATA_W 32
`define IOB_UUT_ADDR_W (12+2)
`define IOB_UUT_AXI_ID_W 1
`define IOB_UUT_AXI_ADDR_W 14
`define IOB_UUT_AXI_DATA_W DATA_W
`define IOB_UUT_AXI_LEN_W 8
`define IOB_UUT_PHY_RST_CNT 20'h00100
`define IOB_UUT_BD_NUM_LOG2 7
`define IOB_UUT_BUFFER_W 11
// Core Configuration Macros.
`define IOB_UUT_VERSION 24'h008100
