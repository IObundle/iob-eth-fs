// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_GRAY_COUNTER_W 1
// Core Configuration Macros.
`define IOB_GRAY_COUNTER_VERSION 24'h008100
