// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_DMA_DATA_W 32
`define IOB_DMA_ADDR_W 5
`define IOB_DMA_AXI_ADDR_W 1
`define IOB_DMA_AXI_LEN_W 8
`define IOB_DMA_AXI_DATA_W 32
`define IOB_DMA_AXI_ID_W 1
`define IOB_DMA_WLEN_W 12
`define IOB_DMA_RLEN_W 12
// Core Configuration Macros.
`define IOB_DMA_VERSION 24'h008100
