// general_operation: General operation group
// Core Configuration Macros.
`define IOB_ETH_TX_VERSION 24'h008100
