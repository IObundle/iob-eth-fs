// general_operation: General operation group
// Core Configuration Macros.
`define IOB_RESET_SYNC_VERSION 24'h008100
