// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_RAM_AT2P_DATA_W 32
`define IOB_RAM_AT2P_ADDR_W 1
// Core Configuration Macros.
`define IOB_RAM_AT2P_VERSION 24'h008100
