// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_ETH_LOGIC_BUFFER_W 11
// Core Configuration Macros.
`define IOB_ETH_LOGIC_VERSION 24'h008100
