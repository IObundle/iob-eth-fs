// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXISTREAM_OUT_CSRS_DATA_W 32
`define IOB_AXISTREAM_OUT_CSRS_TDATA_W 8
`define IOB_AXISTREAM_OUT_CSRS_FIFO_ADDR_W 4
// Core Configuration Macros.
`define IOB_AXISTREAM_OUT_CSRS_SOFT_RESET_ADDR 0
`define IOB_AXISTREAM_OUT_CSRS_SOFT_RESET_W 8
`define IOB_AXISTREAM_OUT_CSRS_ENABLE_ADDR 1
`define IOB_AXISTREAM_OUT_CSRS_ENABLE_W 8
`define IOB_AXISTREAM_OUT_CSRS_DATA_ADDR 4
`define IOB_AXISTREAM_OUT_CSRS_DATA_W 32
`define IOB_AXISTREAM_OUT_CSRS_MODE_ADDR 8
`define IOB_AXISTREAM_OUT_CSRS_MODE_W 8
`define IOB_AXISTREAM_OUT_CSRS_NWORDS_ADDR 12
`define IOB_AXISTREAM_OUT_CSRS_NWORDS_W 32
`define IOB_AXISTREAM_OUT_CSRS_FIFO_FULL_ADDR 16
`define IOB_AXISTREAM_OUT_CSRS_FIFO_FULL_W 8
`define IOB_AXISTREAM_OUT_CSRS_FIFO_EMPTY_ADDR 17
`define IOB_AXISTREAM_OUT_CSRS_FIFO_EMPTY_W 8
`define IOB_AXISTREAM_OUT_CSRS_FIFO_THRESHOLD_ADDR 20
`define IOB_AXISTREAM_OUT_CSRS_FIFO_THRESHOLD_W 32
`define IOB_AXISTREAM_OUT_CSRS_FIFO_LEVEL_ADDR 24
`define IOB_AXISTREAM_OUT_CSRS_FIFO_LEVEL_W 32
`define IOB_AXISTREAM_OUT_CSRS_VERSION_ADDR 28
`define IOB_AXISTREAM_OUT_CSRS_VERSION_W 32
`define IOB_AXISTREAM_OUT_CSRS_VERSION 24'h008100
// Core Derived Parameters. DO NOT CHANGE
`define IOB_AXISTREAM_OUT_CSRS_ADDR_W 5
